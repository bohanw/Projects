module input_assumption(output logic ok);
   assign ok=1'b1;
endmodule
